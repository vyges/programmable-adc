//=============================================================================
// Sample & Hold (S/H) Module
//=============================================================================
// Description: Track and Hold circuit using switched capacitor architecture.
//              Hold time > 200 ns, droop rate < 1 LSB/μs, aperture jitter < 1 ps RMS.
//
// Architecture: Switched capacitor track and hold
// Author:       Vyges Development Team
// Created:      2025-01-27
//=============================================================================

module sample_hold (
    // Clock and Reset
    input  wire        clk,            // System clock
    input  wire        reset_n,        // Reset (active low)
    input  wire        enable,         // S/H enable
    
    // Control
    input  wire        sample_en,      // Sample enable (active high)
    
    // Analog Inputs (digital representation for simulation)
    input  wire [15:0] vin_p,          // Positive input
    input  wire [15:0] vin_n,          // Negative input
    
    // Analog Outputs (digital representation for simulation)
    output reg  [15:0] vout_p,         // Positive output
    output reg  [15:0] vout_n          // Negative output
);

    // Internal signals
    reg [15:0] hold_p, hold_n;         // Hold capacitors (simplified)
    reg        track_mode;             // Track mode indicator
    
    // Track/Hold state machine
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            track_mode <= 1'b0;
            hold_p <= 16'h0000;
            hold_n <= 16'h0000;
        end else if (enable) begin
            if (sample_en) begin
                // Track mode - sample input
                track_mode <= 1'b1;
                hold_p <= vin_p;
                hold_n <= vin_n;
            end else begin
                // Hold mode - maintain sampled value
                track_mode <= 1'b0;
                // hold_p and hold_n maintain their values
            end
        end else begin
            track_mode <= 1'b0;
            hold_p <= 16'h0000;
            hold_n <= 16'h0000;
        end
    end
    
    // Output generation
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            vout_p <= 16'h0000;
            vout_n <= 16'h0000;
        end else if (enable) begin
            if (track_mode) begin
                // Track mode - pass through input
                vout_p <= vin_p;
                vout_n <= vin_n;
            end else begin
                // Hold mode - output held value
                vout_p <= hold_p;
                vout_n <= hold_n;
            end
        end else begin
            vout_p <= 16'h0000;
            vout_n <= 16'h0000;
        end
    end

endmodule 