//=============================================================================
// Programmable ADC - SAR DAC Circuit Implementation (Cadence PDK)
//=============================================================================
// Description: SAR DAC array optimized for Cadence PDK
//              Uses behavioral models and specifications from /docs
// Author: Vyges IP Development Team
// Date: 2025
//=============================================================================

`include "disciplines.vams"

module sar_dac_circuit_cadence #(
    parameter int  RESOLUTION = 16,
    parameter real VDDA = 2.8,
    parameter real VDDD = 1.1,
    parameter real VREF = 2.8,
    parameter real CUNIT = 1e-15,
    parameter real CMISMATCH = 0.001,
    parameter real TEMP_COEF = 20e-6,
    parameter real VOLT_COEF = 50e-6,
    parameter real TEMP = 27.0
)(
    // Clock and control
    input  logic        clk_i,
    input  logic        reset_n_i,
    input  logic        enable_i,
    
    // Resolution control
    input  logic [1:0]  resolution_i,
    
    // DAC control
    input  logic [15:0] dac_code_i,
    input  logic        dac_valid_i,
    input  logic        reset_dac_i,
    
    // Calibration control
    input  logic        cal_enable_i,
    input  logic [7:0]  cal_code_i,
    input  logic        cal_valid_i,
    
    // Analog outputs (electrical discipline)
    output electrical   dac_out_p_o,
    output electrical   dac_out_n_o,
    output electrical   dac_cm_o,
    
    // Status and control
    output logic        ready_o,
    output logic        busy_o,
    output real         dnl_o,
    output real         inl_o,
    output real         temp_drift_o,
    output real         voltage_drift_o
);

    //=============================================================================
    // Cadence PDK specific parameters
    //=============================================================================
    
    // Process parameters from Cadence PDK
    parameter real VTN = 0.45;      // NMOS threshold voltage
    parameter real VTP = -0.45;     // PMOS threshold voltage
    parameter real KP_N = 200e-6;   // NMOS transconductance parameter
    parameter real KP_P = 80e-6;    // PMOS transconductance parameter
    parameter real LAMBDA_N = 0.1;  // NMOS channel length modulation
    parameter real LAMBDA_P = 0.1;  // PMOS channel length modulation
    
    // Capacitor parameters from component specifications
    parameter real C_METAL_METAL = 1e-15;  // Metal-metal capacitor density
    parameter real C_POLY_POLY = 1e-15;    // Poly-poly capacitor density
    parameter real C_MOS = 1e-15;          // MOS capacitor density
    
    //=============================================================================
    // Internal signals and parameters
    //=============================================================================
    
    // Resolution-dependent parameters
    int effective_resolution;
    int max_code;
    real lsb_size;
    
    // Capacitor array signals (electrical discipline)
    electrical cap_array [0:15];  // 16-bit capacitor array
    electrical cap_mismatch [0:15];  // Capacitor mismatch errors
    electrical cap_temp_drift [0:15];  // Temperature drift
    electrical cap_voltage_drift [0:15];  // Voltage drift
    
    // Switch control signals
    logic [15:0] switch_high, switch_low, switch_mid;
    logic [15:0] switch_high_d, switch_low_d, switch_mid_d;
    
    // DAC output signals
    electrical dac_voltage_p, dac_voltage_n;
    electrical dac_voltage_diff, dac_voltage_cm;
    
    // Calibration signals
    real cal_offset, cal_gain;
    real cal_temp_coef, cal_voltage_coef;
    logic [7:0] cal_code_sync;
    
    // Performance monitoring
    real dnl_error, inl_error;
    real temp_error, voltage_error;
    
    // Timing signals
    logic settling_done, conversion_done;
    real settling_time, conversion_time;
    
    // Power supply signals
    electrical vdda, vssa, vref;
    
    //=============================================================================
    // Power supply connections
    //=============================================================================
    
    assign vdda = VDDA;
    assign vssa = 0.0;
    assign vref = VREF;
    
    //=============================================================================
    // Resolution and parameter calculation
    //=============================================================================
    
    // Resolution calculation
    always_comb begin
        case (resolution_i)
            2'b00: effective_resolution = 12;
            2'b01: effective_resolution = 14;
            2'b10: effective_resolution = 16;
            default: effective_resolution = 16;
        endcase
        
        max_code = (1 << effective_resolution) - 1;
        lsb_size = VREF / (1 << effective_resolution);
    end
    
    //=============================================================================
    // Capacitor array initialization (Cadence behavioral)
    //=============================================================================
    
    // Capacitor array generation using Cadence behavioral models
    genvar i;
    generate
        for (i = 0; i < 16; i = i + 1) begin : cap_array_gen
            // Binary-weighted capacitor values
            analog begin
                if (i < effective_resolution) begin
                    // Capacitor value calculation
                    real cap_value = CUNIT * (1 << i);
                    
                    // Capacitor mismatch modeling from component specs
                    real mismatch_factor = 1.0 + CMISMATCH * ($random() - 0.5);
                    real cap_mismatch_value = cap_value * (mismatch_factor - 1.0);
                    
                    // Temperature drift modeling
                    real temp_change = TEMP - 27.0;  // Temperature change from nominal
                    real cap_temp_drift_value = cap_value * TEMP_COEF * temp_change;
                    
                    // Voltage drift modeling
                    real voltage_change = V(vref) - 2.8;  // Voltage change from nominal
                    real cap_voltage_drift_value = cap_value * VOLT_COEF * voltage_change;
                    
                    // Total capacitor value with all effects
                    real total_cap_value = cap_value + cap_mismatch_value + 
                                         cap_temp_drift_value + cap_voltage_drift_value;
                    
                    // Capacitor behavioral model
                    I(cap_array[i]) <+ ddt(total_cap_value * V(cap_array[i]));
                    
                    // Mismatch and drift monitoring
                    V(cap_mismatch[i]) <+ cap_mismatch_value;
                    V(cap_temp_drift[i]) <+ cap_temp_drift_value;
                    V(cap_voltage_drift[i]) <+ cap_voltage_drift_value;
                end else begin
                    // Unused capacitors
                    I(cap_array[i]) <+ 0.0;
                    V(cap_mismatch[i]) <+ 0.0;
                    V(cap_temp_drift[i]) <+ 0.0;
                    V(cap_voltage_drift[i]) <+ 0.0;
                end
            end
        end
    endgenerate
    
    //=============================================================================
    // Switch control logic
    //=============================================================================
    
    // Switch control generation
    always_comb begin
        for (int i = 0; i < 16; i = i + 1) begin
            if (i < effective_resolution) begin
                // DAC code bit determines switch position
                switch_high[i] = dac_code_i[i] && !reset_dac_i;
                switch_low[i] = !dac_code_i[i] && !reset_dac_i;
                switch_mid[i] = reset_dac_i;  // Midscale reset
            end else begin
                // Unused capacitors connected to midscale
                switch_high[i] = 1'b0;
                switch_low[i] = 1'b0;
                switch_mid[i] = 1'b1;
            end
        end
    end
    
    // Synchronize switch signals
    always_ff @(posedge clk_i or negedge reset_n_i) begin
        if (!reset_n_i) begin
            switch_high_d <= 16'h0000;
            switch_low_d <= 16'h0000;
            switch_mid_d <= 16'h0000;
        end else begin
            switch_high_d <= switch_high;
            switch_low_d <= switch_low;
            switch_mid_d <= switch_mid;
        end
    end
    
    //=============================================================================
    // DAC voltage calculation (Cadence behavioral)
    //=============================================================================
    
    // DAC output voltage calculation using Cadence behavioral models
    analog begin
        real total_cap_high = 0.0;
        real total_cap_low = 0.0;
        real total_cap_mid = 0.0;
        real total_cap = 0.0;
        
        // Calculate total capacitance for each switch position
        for (int i = 0; i < 16; i = i + 1) begin
            real cap_value = CUNIT * (1 << i);
            real cap_mismatch_value = V(cap_mismatch[i]);
            real cap_temp_drift_value = V(cap_temp_drift[i]);
            real cap_voltage_drift_value = V(cap_voltage_drift[i]);
            
            real total_cap_value = cap_value + cap_mismatch_value + 
                                 cap_temp_drift_value + cap_voltage_drift_value;
            
            if (switch_high_d[i]) begin
                total_cap_high = total_cap_high + total_cap_value;
            end else if (switch_low_d[i]) begin
                total_cap_low = total_cap_low + total_cap_value;
            end else if (switch_mid_d[i]) begin
                total_cap_mid = total_cap_mid + total_cap_value;
            end
            
            total_cap = total_cap + total_cap_value;
        end
        
        // DAC voltage calculation using charge conservation
        real vhigh = V(vref);
        real vlow = 0.0;
        real vmid = V(vref) / 2.0;
        
        // Charge conservation: Q = C * V
        real total_charge = total_cap_high * vhigh + 
                          total_cap_low * vlow + 
                          total_cap_mid * vmid;
        
        V(dac_voltage_cm) <+ total_charge / total_cap;
        
        // Differential output calculation
        real ideal_voltage = (dac_code_i * V(vref)) / (1 << effective_resolution);
        real voltage_error = V(dac_voltage_cm) - ideal_voltage;
        
        // Apply calibration
        V(dac_voltage_p) <+ V(dac_voltage_cm) + cal_offset + cal_gain * voltage_error;
        V(dac_voltage_n) <+ V(vref) - V(dac_voltage_p);
        V(dac_voltage_diff) <+ V(dac_voltage_p) - V(dac_voltage_n);
        
        // Output assignment
        V(dac_out_p_o) <+ V(dac_voltage_p);
        V(dac_out_n_o) <+ V(dac_voltage_n);
        V(dac_cm_o) <+ V(dac_voltage_cm);
    end
    
    //=============================================================================
    // Calibration implementation
    //=============================================================================
    
    // Calibration code synchronization
    always_ff @(posedge clk_i or negedge reset_n_i) begin
        if (!reset_n_i) begin
            cal_code_sync <= 8'h00;
        end else if (cal_valid_i) begin
            cal_code_sync <= cal_code_i;
        end
    end
    
    // Calibration parameter calculation
    always_comb begin
        if (cal_enable_i) begin
            // Calibration offset (8-bit resolution)
            cal_offset = (cal_code_sync[3:0] - 8.0) * lsb_size / 16.0;
            
            // Calibration gain (8-bit resolution)
            cal_gain = 1.0 + (cal_code_sync[7:4] - 8.0) * 0.001;  // ±0.5% gain adjustment
            
            // Temperature coefficient calibration
            cal_temp_coef = TEMP_COEF * (1.0 + (cal_code_sync[5:4] - 2.0) * 0.1);
            
            // Voltage coefficient calibration
            cal_voltage_coef = VOLT_COEF * (1.0 + (cal_code_sync[7:6] - 2.0) * 0.1);
        end else begin
            cal_offset = 0.0;
            cal_gain = 1.0;
            cal_temp_coef = TEMP_COEF;
            cal_voltage_coef = VOLT_COEF;
        end
    end
    
    //=============================================================================
    // Performance measurement (Cadence behavioral)
    //=============================================================================
    
    // DNL calculation
    analog begin
        real ideal_step = lsb_size;
        real actual_step = V(dac_voltage_diff) / max_code;
        dnl_error = (actual_step - ideal_step) / ideal_step;
    end
    
    // INL calculation
    analog begin
        real ideal_voltage = (dac_code_i * V(vref)) / (1 << effective_resolution);
        real actual_voltage = V(dac_voltage_cm);
        inl_error = (actual_voltage - ideal_voltage) / lsb_size;
    end
    
    // Temperature drift calculation
    analog begin
        real temp_change = TEMP - 27.0;  // Temperature change from nominal
        temp_error = temp_change * cal_temp_coef;
    end
    
    // Voltage drift calculation
    analog begin
        real voltage_change = V(vref) - 2.8;  // Voltage change from nominal
        voltage_error = voltage_change * cal_voltage_coef;
    end
    
    //=============================================================================
    // Timing and control logic
    //=============================================================================
    
    // Settling time calculation
    analog begin
        real total_cap = 0.0;
        real switch_resistance = 200.0;  // 200Ω switch resistance from specs
        
        for (int i = 0; i < 16; i = i + 1) begin
            total_cap = total_cap + CUNIT * (1 << i);
        end
        
        real tau = switch_resistance * total_cap;
        settling_time = 5.0 * tau;  // 5 time constants for settling
    end
    
    // Conversion timing
    always_ff @(posedge clk_i or negedge reset_n_i) begin
        if (!reset_n_i) begin
            settling_done <= 1'b0;
            conversion_done <= 1'b0;
            conversion_time <= 0.0;
        end else begin
            if (dac_valid_i) begin
                settling_done <= 1'b0;
                conversion_done <= 1'b0;
                conversion_time <= 0.0;
            end else begin
                conversion_time <= conversion_time + 10e-9;  // 10ns increment
                
                if (conversion_time >= settling_time) begin
                    settling_done <= 1'b1;
                end
                
                if (conversion_time >= settling_time + 100e-9) begin
                    conversion_done <= 1'b1;
                end
            end
        end
    end
    
    // Ready and busy signals
    always_ff @(posedge clk_i or negedge reset_n_i) begin
        if (!reset_n_i) begin
            ready_o <= 1'b0;
            busy_o <= 1'b0;
        end else begin
            ready_o <= enable_i && !dac_valid_i;
            busy_o <= dac_valid_i || !settling_done;
        end
    end
    
    //=============================================================================
    // Output assignment
    //=============================================================================
    
    // Performance output assignment
    always_comb begin
        dnl_o = dnl_error;
        inl_o = inl_error;
        temp_drift_o = temp_error;
        voltage_drift_o = voltage_error;
    end
    
    //=============================================================================
    // Power consumption calculation (Cadence behavioral)
    //=============================================================================
    
    // Static power calculation
    analog begin
        real leakage_current = 10e-9;  // 10nA leakage current from specs
        real static_power = leakage_current * V(vdda);
        
        // Dynamic power calculation
        real switching_freq = 5e6;    // 5MHz switching frequency
        real total_cap = 0.0;
        
        for (int i = 0; i < 16; i = i + 1) begin
            total_cap = total_cap + CUNIT * (1 << i);
        end
        
        real dynamic_power = 0.5 * total_cap * V(vdda) * V(vdda) * switching_freq;
        
        // Total power monitoring
        real total_power = static_power + dynamic_power;
    end
    
    //=============================================================================
    // Cadence-specific assertions and coverage
    //=============================================================================
    
    // Input range assertion
    property input_range_check;
        @(posedge clk_i) disable iff (!reset_n_i)
        (dac_code_i >= 0) && (dac_code_i <= max_code);
    endproperty
    
    assert property (input_range_check)
    else $error("DAC input code out of range");
    
    // Output range assertion
    property output_range_check;
        @(posedge clk_i) disable iff (!reset_n_i)
        (V(dac_out_p_o) >= 0) && (V(dac_out_p_o) <= VREF) &&
        (V(dac_out_n_o) >= 0) && (V(dac_out_n_o) <= VREF);
    endproperty
    
    assert property (output_range_check)
    else $error("DAC output voltage out of range");
    
    // Resolution coverage
    covergroup resolution_coverage @(posedge clk_i);
        resolution_cp: coverpoint resolution_i {
            bins res_12bit = {2'b00};
            bins res_14bit = {2'b01};
            bins res_16bit = {2'b10};
            bins invalid = {2'b11};
        }
    endgroup
    
    resolution_coverage res_cov = new();
    
    //=============================================================================
    // Cadence-specific performance monitoring
    //=============================================================================
    
    // DNL monitoring
    always @(posedge clk_i) begin
        if (conversion_done) begin
            if (abs(dnl_error) > 0.5) begin
                $warning("DAC DNL error: %f LSB", dnl_error);
            end
        end
    end
    
    // INL monitoring
    always @(posedge clk_i) begin
        if (conversion_done) begin
            if (abs(inl_error) > 1.0) begin
                $warning("DAC INL error: %f LSB", inl_error);
            end
        end
    end
    
    // Temperature drift monitoring
    always @(posedge clk_i) begin
        if (conversion_done) begin
            if (abs(temp_error) > 1e-3) begin
                $warning("DAC temperature drift: %f V", temp_error);
            end
        end
    end
    
endmodule 