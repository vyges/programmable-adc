//=============================================================================
// SAR Controller Module
//=============================================================================
// Description: Successive Approximation Register controller for ADC conversion.
//              Supports 12, 14, 16-bit resolution with configurable conversion time.
//              Conversion time: 200 ns (5 MSPS), power < 3 mW.
//
// Architecture: Successive Approximation
// Author:       Vyges Development Team
// Created:      2025-01-27
//=============================================================================

module sar_controller (
    // Clock and Reset
    input  wire        clk,            // System clock
    input  wire        reset_n,        // Reset (active low)
    input  wire        enable,         // SAR enable
    
    // Control
    input  wire        start_conv,     // Start conversion
    input  wire [1:0]  resolution,     // Resolution (00=12bit, 01=14bit, 10=16bit)
    input  wire        auto_mode,      // Auto conversion mode
    
    // Analog Inputs (digital representation for simulation)
    input  wire [15:0] vin_p,          // Positive input
    input  wire [15:0] vin_n,          // Negative input
    
    // DAC Interface
    output reg  [15:0] dac_out_p,      // DAC positive output
    output reg  [15:0] dac_out_n,      // DAC negative output
    input  wire        comp_out,       // Comparator output
    
    // Output
    output reg  [15:0] data_out,       // Conversion result
    output reg         busy,           // Conversion busy
    output reg         valid           // Data valid
);

    // State machine states
    localparam IDLE = 3'b000;
    localparam SAMPLE = 3'b001;
    localparam CONVERT = 3'b010;
    localparam DONE = 3'b011;
    
    reg [2:0] state, next_state;
    reg [4:0] bit_counter;             // Bit counter for conversion
    reg [15:0] sar_register;           // SAR register
    reg [15:0] max_bits;               // Maximum bits based on resolution
    
    // State machine
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            state <= IDLE;
        end else begin
            state <= next_state;
        end
    end
    
    // Next state logic
    always @(*) begin
        case (state)
            IDLE: begin
                if (start_conv && enable) begin
                    next_state = SAMPLE;
                end else begin
                    next_state = IDLE;
                end
            end
            
            SAMPLE: begin
                next_state = CONVERT;
            end
            
            CONVERT: begin
                if (bit_counter == 5'h0) begin
                    next_state = DONE;
                end else begin
                    next_state = CONVERT;
                end
            end
            
            DONE: begin
                if (auto_mode && enable) begin
                    next_state = SAMPLE;
                end else begin
                    next_state = IDLE;
                end
            end
            
            default: next_state = IDLE;
        endcase
    end
    
    // Resolution setting
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            max_bits <= 16'h0010;  // Default 16-bit
        end else begin
            case (resolution)
                2'b00: max_bits <= 16'h000C;  // 12-bit
                2'b01: max_bits <= 16'h000E;  // 14-bit
                2'b10: max_bits <= 16'h0010;  // 16-bit
                default: max_bits <= 16'h0010;
            endcase
        end
    end
    
    // Bit counter and SAR logic
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            bit_counter <= 5'h0;
            sar_register <= 16'h0000;
            busy <= 1'b0;
            valid <= 1'b0;
            data_out <= 16'h0000;
        end else begin
            case (state)
                IDLE: begin
                    busy <= 1'b0;
                    valid <= 1'b0;
                    bit_counter <= 5'h0;
                    sar_register <= 16'h0000;
                end
                
                SAMPLE: begin
                    busy <= 1'b1;
                    valid <= 1'b0;
                    bit_counter <= max_bits[4:0] - 1;  // Start from MSB
                    sar_register <= 16'h0000;
                end
                
                CONVERT: begin
                    busy <= 1'b1;
                    valid <= 1'b0;
                    
                    if (comp_out) begin
                        // Input > DAC, set current bit
                        sar_register[bit_counter] <= 1'b1;
                    end else begin
                        // Input <= DAC, clear current bit
                        sar_register[bit_counter] <= 1'b0;
                    end
                    
                    if (bit_counter > 0) begin
                        bit_counter <= bit_counter - 1;
                    end
                end
                
                DONE: begin
                    busy <= 1'b0;
                    valid <= 1'b1;
                    data_out <= sar_register;
                end
                
                default: begin
                    busy <= 1'b0;
                    valid <= 1'b0;
                end
            endcase
        end
    end
    
    // DAC output generation based on SAR register
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            dac_out_p <= 16'h0000;
            dac_out_n <= 16'h0000;
        end else if (state == CONVERT) begin
            // Generate DAC output based on current SAR register value
            // This is a simplified representation for simulation
            dac_out_p <= sar_register;
            dac_out_n <= 16'h0000;
        end else begin
            dac_out_p <= 16'h0000;
            dac_out_n <= 16'h0000;
        end
    end

endmodule 